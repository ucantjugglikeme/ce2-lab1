module smooth_sorter#(
    parameter n = 256
)(
    input clk,
    input [31:0] dataIn,
    input is_input,
    input i,
    output [31:0] dataOut
);



endmodule
